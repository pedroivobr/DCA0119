library verilog;
use verilog.vl_types.all;
entity main_vlg_check_tst is
    port(
        resultado       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end main_vlg_check_tst;
