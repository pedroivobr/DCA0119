library verilog;
use verilog.vl_types.all;
entity timeSelector_vlg_vec_tst is
end timeSelector_vlg_vec_tst;
