library verilog;
use verilog.vl_types.all;
entity testes_vlg_check_tst is
    port(
        pin_name2       : in     vl_logic;
        pin_name3       : in     vl_logic;
        pin_name4       : in     vl_logic;
        pin_name5       : in     vl_logic;
        pin_name6       : in     vl_logic;
        pin_name7       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end testes_vlg_check_tst;
