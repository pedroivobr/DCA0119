-- megafunction wizard: %ALTFP_CONVERT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_CONVERT 

-- ============================================================
-- File Name: altfp_convert1.vhd
-- Megafunction Name(s):
-- 			ALTFP_CONVERT
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altfp_convert CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" OPERATION="FLOAT2INT" ROUNDING="TO_NEAREST" WIDTH_DATA=32 WIDTH_EXP_INPUT=8 WIDTH_EXP_OUTPUT=8 WIDTH_INT=32 WIDTH_MAN_INPUT=23 WIDTH_MAN_OUTPUT=23 WIDTH_RESULT=32 clock dataa result
--VERSION_BEGIN 13.0 cbx_altbarrel_shift 2013:06:12:18:03:43:SJ cbx_altfp_convert 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_altsyncram 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_abs 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_lpm_decode 2013:06:12:18:03:43:SJ cbx_lpm_divide 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_stratixiii 2013:06:12:18:03:43:SJ cbx_stratixv 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" PIPELINE=2 SHIFTDIR="LEFT" SHIFTTYPE="LOGICAL" WIDTH=54 WIDTHDIST=6 aclr clk_en clock data distance result
--VERSION_BEGIN 13.0 cbx_altbarrel_shift 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = reg 113 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert1_altbarrel_shift_grf IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (53 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (5 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (53 DOWNTO 0)
	 ); 
 END altfp_convert1_altbarrel_shift_grf;

 ARCHITECTURE RTL OF altfp_convert1_altbarrel_shift_grf IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(53 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper2d	:	STD_LOGIC_VECTOR(53 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec3r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec4r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec5r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range287w300w301w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range287w296w297w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range308w321w322w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range308w317w318w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range330w343w344w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range330w339w340w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range353w365w366w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range353w361w362w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range372w384w385w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range372w380w381w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range393w405w406w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range393w401w402w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range287w292w293w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range308w313w314w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range330w335w336w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range353w357w358w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range372w376w377w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range393w397w398w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range287w300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range287w296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range308w321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range308w317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range330w343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range330w339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range353w365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range353w361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range372w384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range372w380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range393w405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range393w401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_dir_w_range284w299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_dir_w_range306w320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_dir_w_range327w342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_dir_w_range351w364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_dir_w_range370w383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_dir_w_range390w404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range287w292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range308w313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range330w335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range353w357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range372w376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range393w397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range287w300w301w302w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range308w321w322w323w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range330w343w344w345w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range353w365w366w367w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range372w384w385w386w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range393w405w406w407w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w303w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w324w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w346w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w368w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w387w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w408w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (377 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (323 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w295w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w298w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w316w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w319w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w338w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w341w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w360w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w363w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w379w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w382w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w400w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w403w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_dir_w_range284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_dir_w_range306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_dir_w_range327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_dir_w_range351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_dir_w_range370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_dir_w_range390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sbit_w_range305w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sbit_w_range325w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sbit_w_range347w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sbit_w_range369w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sbit_w_range388w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sbit_w_range282w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sel_w_range287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sel_w_range308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sel_w_range330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sel_w_range353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sel_w_range372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sel_w_range393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_smux_w_range334w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_smux_w_range396w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range287w300w301w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range287w300w(0) AND wire_altbarrel_shift6_w298w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range287w296w297w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range287w296w(0) AND wire_altbarrel_shift6_w295w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range308w321w322w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range308w321w(0) AND wire_altbarrel_shift6_w319w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range308w317w318w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range308w317w(0) AND wire_altbarrel_shift6_w316w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range330w343w344w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range330w343w(0) AND wire_altbarrel_shift6_w341w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range330w339w340w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range330w339w(0) AND wire_altbarrel_shift6_w338w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range353w365w366w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range353w365w(0) AND wire_altbarrel_shift6_w363w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range353w361w362w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range353w361w(0) AND wire_altbarrel_shift6_w360w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range372w384w385w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range372w384w(0) AND wire_altbarrel_shift6_w382w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range372w380w381w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range372w380w(0) AND wire_altbarrel_shift6_w379w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range393w405w406w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range393w405w(0) AND wire_altbarrel_shift6_w403w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range393w401w402w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range393w401w(0) AND wire_altbarrel_shift6_w400w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range287w292w293w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range287w292w(0) AND wire_altbarrel_shift6_w_sbit_w_range282w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range308w313w314w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range308w313w(0) AND wire_altbarrel_shift6_w_sbit_w_range305w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range330w335w336w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range330w335w(0) AND wire_altbarrel_shift6_w_sbit_w_range325w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range353w357w358w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range353w357w(0) AND wire_altbarrel_shift6_w_sbit_w_range347w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range372w376w377w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range372w376w(0) AND wire_altbarrel_shift6_w_sbit_w_range369w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range393w397w398w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range393w397w(0) AND wire_altbarrel_shift6_w_sbit_w_range388w(i);
	END GENERATE loop17;
	wire_altbarrel_shift6_w_lg_w_sel_w_range287w300w(0) <= wire_altbarrel_shift6_w_sel_w_range287w(0) AND wire_altbarrel_shift6_w_lg_w_dir_w_range284w299w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range287w296w(0) <= wire_altbarrel_shift6_w_sel_w_range287w(0) AND wire_altbarrel_shift6_w_dir_w_range284w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range308w321w(0) <= wire_altbarrel_shift6_w_sel_w_range308w(0) AND wire_altbarrel_shift6_w_lg_w_dir_w_range306w320w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range308w317w(0) <= wire_altbarrel_shift6_w_sel_w_range308w(0) AND wire_altbarrel_shift6_w_dir_w_range306w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range330w343w(0) <= wire_altbarrel_shift6_w_sel_w_range330w(0) AND wire_altbarrel_shift6_w_lg_w_dir_w_range327w342w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range330w339w(0) <= wire_altbarrel_shift6_w_sel_w_range330w(0) AND wire_altbarrel_shift6_w_dir_w_range327w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range353w365w(0) <= wire_altbarrel_shift6_w_sel_w_range353w(0) AND wire_altbarrel_shift6_w_lg_w_dir_w_range351w364w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range353w361w(0) <= wire_altbarrel_shift6_w_sel_w_range353w(0) AND wire_altbarrel_shift6_w_dir_w_range351w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range372w384w(0) <= wire_altbarrel_shift6_w_sel_w_range372w(0) AND wire_altbarrel_shift6_w_lg_w_dir_w_range370w383w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range372w380w(0) <= wire_altbarrel_shift6_w_sel_w_range372w(0) AND wire_altbarrel_shift6_w_dir_w_range370w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range393w405w(0) <= wire_altbarrel_shift6_w_sel_w_range393w(0) AND wire_altbarrel_shift6_w_lg_w_dir_w_range390w404w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range393w401w(0) <= wire_altbarrel_shift6_w_sel_w_range393w(0) AND wire_altbarrel_shift6_w_dir_w_range390w(0);
	wire_altbarrel_shift6_w_lg_w_dir_w_range284w299w(0) <= NOT wire_altbarrel_shift6_w_dir_w_range284w(0);
	wire_altbarrel_shift6_w_lg_w_dir_w_range306w320w(0) <= NOT wire_altbarrel_shift6_w_dir_w_range306w(0);
	wire_altbarrel_shift6_w_lg_w_dir_w_range327w342w(0) <= NOT wire_altbarrel_shift6_w_dir_w_range327w(0);
	wire_altbarrel_shift6_w_lg_w_dir_w_range351w364w(0) <= NOT wire_altbarrel_shift6_w_dir_w_range351w(0);
	wire_altbarrel_shift6_w_lg_w_dir_w_range370w383w(0) <= NOT wire_altbarrel_shift6_w_dir_w_range370w(0);
	wire_altbarrel_shift6_w_lg_w_dir_w_range390w404w(0) <= NOT wire_altbarrel_shift6_w_dir_w_range390w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range287w292w(0) <= NOT wire_altbarrel_shift6_w_sel_w_range287w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range308w313w(0) <= NOT wire_altbarrel_shift6_w_sel_w_range308w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range330w335w(0) <= NOT wire_altbarrel_shift6_w_sel_w_range330w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range353w357w(0) <= NOT wire_altbarrel_shift6_w_sel_w_range353w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range372w376w(0) <= NOT wire_altbarrel_shift6_w_sel_w_range372w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range393w397w(0) <= NOT wire_altbarrel_shift6_w_sel_w_range393w(0);
	loop18 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range287w300w301w302w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range287w300w301w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range287w296w297w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range308w321w322w323w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range308w321w322w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range308w317w318w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range330w343w344w345w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range330w343w344w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range330w339w340w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range353w365w366w367w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range353w365w366w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range353w361w362w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range372w384w385w386w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range372w384w385w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range372w380w381w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range393w405w406w407w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range393w405w406w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range393w401w402w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w303w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range287w300w301w302w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range287w292w293w(i);
	END GENERATE loop24;
	loop25 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w324w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range308w321w322w323w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range308w313w314w(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w346w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range330w343w344w345w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range330w335w336w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w368w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range353w365w366w367w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range353w357w358w(i);
	END GENERATE loop27;
	loop28 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w387w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range372w384w385w386w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range372w376w377w(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 53 GENERATE 
		wire_altbarrel_shift6_w408w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range393w405w406w407w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range393w397w398w(i);
	END GENERATE loop29;
	dir_w <= ( dir_pipe(1) & dir_w(4 DOWNTO 3) & dir_pipe(0) & dir_w(1 DOWNTO 0) & direction_w);
	direction_w <= '0';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(377 DOWNTO 324);
	sbit_w <= ( sbit_piper2d & smux_w(269 DOWNTO 162) & sbit_piper1d & smux_w(107 DOWNTO 0) & data);
	sel_w <= ( sel_pipec5r1d & sel_pipec4r1d & sel_pipec3r1d & distance(2 DOWNTO 0));
	smux_w <= ( wire_altbarrel_shift6_w408w & wire_altbarrel_shift6_w387w & wire_altbarrel_shift6_w368w & wire_altbarrel_shift6_w346w & wire_altbarrel_shift6_w324w & wire_altbarrel_shift6_w303w);
	wire_altbarrel_shift6_w295w <= ( pad_w(0) & sbit_w(53 DOWNTO 1));
	wire_altbarrel_shift6_w298w <= ( sbit_w(52 DOWNTO 0) & pad_w(0));
	wire_altbarrel_shift6_w316w <= ( pad_w(1 DOWNTO 0) & sbit_w(107 DOWNTO 56));
	wire_altbarrel_shift6_w319w <= ( sbit_w(105 DOWNTO 54) & pad_w(1 DOWNTO 0));
	wire_altbarrel_shift6_w338w <= ( pad_w(3 DOWNTO 0) & sbit_w(161 DOWNTO 112));
	wire_altbarrel_shift6_w341w <= ( sbit_w(157 DOWNTO 108) & pad_w(3 DOWNTO 0));
	wire_altbarrel_shift6_w360w <= ( pad_w(7 DOWNTO 0) & sbit_w(215 DOWNTO 170));
	wire_altbarrel_shift6_w363w <= ( sbit_w(207 DOWNTO 162) & pad_w(7 DOWNTO 0));
	wire_altbarrel_shift6_w379w <= ( pad_w(15 DOWNTO 0) & sbit_w(269 DOWNTO 232));
	wire_altbarrel_shift6_w382w <= ( sbit_w(253 DOWNTO 216) & pad_w(15 DOWNTO 0));
	wire_altbarrel_shift6_w400w <= ( pad_w(31 DOWNTO 0) & sbit_w(323 DOWNTO 302));
	wire_altbarrel_shift6_w403w <= ( sbit_w(291 DOWNTO 270) & pad_w(31 DOWNTO 0));
	wire_altbarrel_shift6_w_dir_w_range284w(0) <= dir_w(0);
	wire_altbarrel_shift6_w_dir_w_range306w(0) <= dir_w(1);
	wire_altbarrel_shift6_w_dir_w_range327w(0) <= dir_w(2);
	wire_altbarrel_shift6_w_dir_w_range351w(0) <= dir_w(3);
	wire_altbarrel_shift6_w_dir_w_range370w(0) <= dir_w(4);
	wire_altbarrel_shift6_w_dir_w_range390w(0) <= dir_w(5);
	wire_altbarrel_shift6_w_sbit_w_range305w <= sbit_w(107 DOWNTO 54);
	wire_altbarrel_shift6_w_sbit_w_range325w <= sbit_w(161 DOWNTO 108);
	wire_altbarrel_shift6_w_sbit_w_range347w <= sbit_w(215 DOWNTO 162);
	wire_altbarrel_shift6_w_sbit_w_range369w <= sbit_w(269 DOWNTO 216);
	wire_altbarrel_shift6_w_sbit_w_range388w <= sbit_w(323 DOWNTO 270);
	wire_altbarrel_shift6_w_sbit_w_range282w <= sbit_w(53 DOWNTO 0);
	wire_altbarrel_shift6_w_sel_w_range287w(0) <= sel_w(0);
	wire_altbarrel_shift6_w_sel_w_range308w(0) <= sel_w(1);
	wire_altbarrel_shift6_w_sel_w_range330w(0) <= sel_w(2);
	wire_altbarrel_shift6_w_sel_w_range353w(0) <= sel_w(3);
	wire_altbarrel_shift6_w_sel_w_range372w(0) <= sel_w(4);
	wire_altbarrel_shift6_w_sel_w_range393w(0) <= sel_w(5);
	wire_altbarrel_shift6_w_smux_w_range334w <= smux_w(161 DOWNTO 108);
	wire_altbarrel_shift6_w_smux_w_range396w <= smux_w(323 DOWNTO 270);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe <= ( dir_w(5) & dir_w(2));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_altbarrel_shift6_w_smux_w_range334w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper2d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper2d <= wire_altbarrel_shift6_w_smux_w_range396w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec3r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec3r1d <= distance(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec4r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec4r1d <= distance(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec5r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec5r1d <= distance(5);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --altfp_convert1_altbarrel_shift_grf

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 5 lpm_compare 4 reg 281 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert1_altfp_convert_3tm IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END altfp_convert1_altfp_convert_3tm;

 ARCHITECTURE RTL OF altfp_convert1_altfp_convert_3tm IS

	 SIGNAL  wire_altbarrel_shift6_result	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL	 added_power2_reg	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit1_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit1_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit1_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit2_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit2_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit2_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_below_lower_limit2_reg3_w_lg_q229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 below_lower_limit2_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_below_lower_limit2_reg4_w_lg_q260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dataa_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 equal_upper_limit_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 equal_upper_limit_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 equal_upper_limit_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_equal_upper_limit_reg3_w_lg_q220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exceed_upper_limit_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exceed_upper_limit_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exceed_upper_limit_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exceed_upper_limit_reg3_w_lg_q221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exceed_upper_limit_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_or_reg4_w_lg_q118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 int_or1_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 int_or2_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 int_or_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 int_or_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_int_or_reg3_w_lg_q219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 integer_result_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 integer_rounded_reg	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lowest_int_sel_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_lowest_int_sel_reg_w_lg_q257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 man_or1_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or2_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_or_reg4_w_lg_q120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 mantissa_input_reg	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 max_shift_exceeder_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 max_shift_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 power2_value_reg	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_input_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_input_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_input_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_sign_input_reg3_w_lg_q222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sign_input_reg3_w_lg_q224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 sign_input_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_sub4_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub5_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_add_sub5_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_add_sub7_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_sub7_datab	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add_sub7_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add_sub8_w_lg_w_lg_cout233w234w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_add_sub8_w_lg_cout232w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_add_sub8_w_lg_cout233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub8_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_sub8_datab	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_add_sub8_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_add_sub9_datab	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_add_sub9_result	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_cmpr1_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr1_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr2_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr3_alb	:	STD_LOGIC;
	 SIGNAL  wire_max_shift_compare_agb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_guard_bit_w201w202w203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_add_1_w206w207w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_below_limit_exceeders267w268w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exceed_limit_exceeders278w279w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_guard_bit_w201w202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_lowest_integer_selector213w214w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sign_input_w238w271w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sign_input_w238w239w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_add_1_w205w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_below_limit_exceeders266w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_exceed_limit_exceeders277w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_lowest_integer_selector212w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_input_w270w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_input_w237w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range8w14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range13w19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range18w24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range23w29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range28w34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range33w39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range38w44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_add_1_w206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_below_limit_exceeders267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_denormal_input_w258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exceed_limit_exceeders278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_guard_bit_w201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_lowest_integer_selector213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_nan_input_w273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_input_w238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_zero_input_w259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_infinity_input_w274w275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_infinity_input_w274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range6w12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range11w17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range16w22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range21w27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range26w32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range31w37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range36w42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range47w51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range74w78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range71w75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range68w72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range65w69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range62w66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range59w63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range56w60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range53w57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range50w54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range84w88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range81w85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range111w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range108w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range105w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range102w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range99w103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range96w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range93w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range90w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range87w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range135w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range165w169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range168w172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range171w175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range174w178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range177w181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range180w184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range183w187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range186w190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range189w193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range192w196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range138w142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range195w199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range141w145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range144w148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range147w151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range150w154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range153w157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range156w160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range159w163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range162w166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  add_1_cout_w :	STD_LOGIC;
	 SIGNAL  add_1_w :	STD_LOGIC;
	 SIGNAL  all_zeroes_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  barrel_mantissa_input :	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  barrel_zero_padding_w :	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  below_limit_exceeders :	STD_LOGIC;
	 SIGNAL  below_limit_integer :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  below_lower_limit1_w :	STD_LOGIC;
	 SIGNAL  below_lower_limit2_w :	STD_LOGIC;
	 SIGNAL  bias_value_less_1_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  bias_value_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  const_bias_value_add_width_res_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  denormal_input_w :	STD_LOGIC;
	 SIGNAL  equal_upper_limit_w :	STD_LOGIC;
	 SIGNAL  exceed_limit_exceeders :	STD_LOGIC;
	 SIGNAL  exceed_limit_integer :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  exceed_upper_limit_w :	STD_LOGIC;
	 SIGNAL  exp_and :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_and_w :	STD_LOGIC;
	 SIGNAL  exp_bus :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_or :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_or_w :	STD_LOGIC;
	 SIGNAL  exponent_input :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  guard_bit_w :	STD_LOGIC;
	 SIGNAL  implied_mantissa_input :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  infinity_input_w :	STD_LOGIC;
	 SIGNAL  infinity_value_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  int_or1_w :	STD_LOGIC;
	 SIGNAL  int_or2_w :	STD_LOGIC;
	 SIGNAL  integer_output :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  integer_post_round :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  integer_pre_round :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  integer_result :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  integer_rounded :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  integer_rounded_tmp :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  integer_tmp_output :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  inv_add_1_adder1_w :	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  inv_add_1_adder2_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  inv_integer :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  lbarrel_shift_result_w :	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  lbarrel_shift_w :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  lower_limit_selector :	STD_LOGIC;
	 SIGNAL  lowest_integer_selector :	STD_LOGIC;
	 SIGNAL  lowest_integer_value :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  man_bus1 :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  man_bus2 :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  man_or1 :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  man_or1_w :	STD_LOGIC;
	 SIGNAL  man_or2 :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  man_or2_w :	STD_LOGIC;
	 SIGNAL  man_or_w :	STD_LOGIC;
	 SIGNAL  mantissa_input :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  max_shift_reg_w :	STD_LOGIC;
	 SIGNAL  max_shift_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  more_than_max_shift_w :	STD_LOGIC;
	 SIGNAL  nan_input_w :	STD_LOGIC;
	 SIGNAL  neg_infi_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  padded_exponent_input :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  pos_infi_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  power2_value_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  round_bit_w :	STD_LOGIC;
	 SIGNAL  sign_input :	STD_LOGIC;
	 SIGNAL  sign_input_w :	STD_LOGIC;
	 SIGNAL  signed_integer :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  sticky_bit_w :	STD_LOGIC;
	 SIGNAL  sticky_bus :	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  sticky_or :	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  unsigned_integer :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  upper_limit_w :	STD_LOGIC;
	 SIGNAL  zero_input_w :	STD_LOGIC;
	 SIGNAL  wire_w_exp_and_range8w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_inv_integer_range218w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  altfp_convert1_altbarrel_shift_grf
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(53 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(53 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_guard_bit_w201w202w203w(0) <= wire_w_lg_w_lg_guard_bit_w201w202w(0) AND sticky_bit_w;
	loop30 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_w_lg_add_1_w206w207w(i) <= wire_w_lg_add_1_w206w(0) AND integer_pre_round(i);
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_lg_below_limit_exceeders267w268w(i) <= wire_w_lg_below_limit_exceeders267w(0) AND integer_output(i);
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_lg_exceed_limit_exceeders278w279w(i) <= wire_w_lg_exceed_limit_exceeders278w(0) AND below_limit_integer(i);
	END GENERATE loop32;
	wire_w_lg_w_lg_guard_bit_w201w202w(0) <= wire_w_lg_guard_bit_w201w(0) AND round_bit_w;
	loop33 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_w_lg_lowest_integer_selector213w214w(i) <= wire_w_lg_lowest_integer_selector213w(0) AND integer_rounded_tmp(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_lg_sign_input_w238w271w(i) <= wire_w_lg_sign_input_w238w(0) AND pos_infi_w(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_w_lg_sign_input_w238w239w(i) <= wire_w_lg_sign_input_w238w(0) AND unsigned_integer(i);
	END GENERATE loop35;
	loop36 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_add_1_w205w(i) <= add_1_w AND integer_post_round(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_below_limit_exceeders266w(i) <= below_limit_exceeders AND all_zeroes_w(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_exceed_limit_exceeders277w(i) <= exceed_limit_exceeders AND infinity_value_w(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_lowest_integer_selector212w(i) <= lowest_integer_selector AND lowest_integer_value(i);
	END GENERATE loop39;
	loop40 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_sign_input_w270w(i) <= sign_input_w AND neg_infi_w(i);
	END GENERATE loop40;
	loop41 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_sign_input_w237w(i) <= sign_input_w AND signed_integer(i);
	END GENERATE loop41;
	wire_w_lg_w_exp_and_range8w14w(0) <= wire_w_exp_and_range8w(0) AND wire_w_exp_bus_range10w(0);
	wire_w_lg_w_exp_and_range13w19w(0) <= wire_w_exp_and_range13w(0) AND wire_w_exp_bus_range15w(0);
	wire_w_lg_w_exp_and_range18w24w(0) <= wire_w_exp_and_range18w(0) AND wire_w_exp_bus_range20w(0);
	wire_w_lg_w_exp_and_range23w29w(0) <= wire_w_exp_and_range23w(0) AND wire_w_exp_bus_range25w(0);
	wire_w_lg_w_exp_and_range28w34w(0) <= wire_w_exp_and_range28w(0) AND wire_w_exp_bus_range30w(0);
	wire_w_lg_w_exp_and_range33w39w(0) <= wire_w_exp_and_range33w(0) AND wire_w_exp_bus_range35w(0);
	wire_w_lg_w_exp_and_range38w44w(0) <= wire_w_exp_and_range38w(0) AND wire_w_exp_bus_range40w(0);
	wire_w_lg_add_1_w206w(0) <= NOT add_1_w;
	wire_w_lg_below_limit_exceeders267w(0) <= NOT below_limit_exceeders;
	wire_w_lg_denormal_input_w258w(0) <= NOT denormal_input_w;
	wire_w_lg_exceed_limit_exceeders278w(0) <= NOT exceed_limit_exceeders;
	wire_w_lg_guard_bit_w201w(0) <= NOT guard_bit_w;
	wire_w_lg_lowest_integer_selector213w(0) <= NOT lowest_integer_selector;
	wire_w_lg_nan_input_w273w(0) <= NOT nan_input_w;
	wire_w_lg_sign_input_w238w(0) <= NOT sign_input_w;
	wire_w_lg_zero_input_w259w(0) <= NOT zero_input_w;
	wire_w_lg_w_lg_infinity_input_w274w275w(0) <= wire_w_lg_infinity_input_w274w(0) OR exceed_upper_limit_reg4;
	wire_w_lg_infinity_input_w274w(0) <= infinity_input_w OR max_shift_exceeder_reg;
	wire_w_lg_w_exp_or_range6w12w(0) <= wire_w_exp_or_range6w(0) OR wire_w_exp_bus_range10w(0);
	wire_w_lg_w_exp_or_range11w17w(0) <= wire_w_exp_or_range11w(0) OR wire_w_exp_bus_range15w(0);
	wire_w_lg_w_exp_or_range16w22w(0) <= wire_w_exp_or_range16w(0) OR wire_w_exp_bus_range20w(0);
	wire_w_lg_w_exp_or_range21w27w(0) <= wire_w_exp_or_range21w(0) OR wire_w_exp_bus_range25w(0);
	wire_w_lg_w_exp_or_range26w32w(0) <= wire_w_exp_or_range26w(0) OR wire_w_exp_bus_range30w(0);
	wire_w_lg_w_exp_or_range31w37w(0) <= wire_w_exp_or_range31w(0) OR wire_w_exp_bus_range35w(0);
	wire_w_lg_w_exp_or_range36w42w(0) <= wire_w_exp_or_range36w(0) OR wire_w_exp_bus_range40w(0);
	wire_w_lg_w_man_or1_range47w51w(0) <= wire_w_man_or1_range47w(0) OR wire_w_man_bus1_range49w(0);
	wire_w_lg_w_man_or1_range74w78w(0) <= wire_w_man_or1_range74w(0) OR wire_w_man_bus1_range76w(0);
	wire_w_lg_w_man_or1_range71w75w(0) <= wire_w_man_or1_range71w(0) OR wire_w_man_bus1_range73w(0);
	wire_w_lg_w_man_or1_range68w72w(0) <= wire_w_man_or1_range68w(0) OR wire_w_man_bus1_range70w(0);
	wire_w_lg_w_man_or1_range65w69w(0) <= wire_w_man_or1_range65w(0) OR wire_w_man_bus1_range67w(0);
	wire_w_lg_w_man_or1_range62w66w(0) <= wire_w_man_or1_range62w(0) OR wire_w_man_bus1_range64w(0);
	wire_w_lg_w_man_or1_range59w63w(0) <= wire_w_man_or1_range59w(0) OR wire_w_man_bus1_range61w(0);
	wire_w_lg_w_man_or1_range56w60w(0) <= wire_w_man_or1_range56w(0) OR wire_w_man_bus1_range58w(0);
	wire_w_lg_w_man_or1_range53w57w(0) <= wire_w_man_or1_range53w(0) OR wire_w_man_bus1_range55w(0);
	wire_w_lg_w_man_or1_range50w54w(0) <= wire_w_man_or1_range50w(0) OR wire_w_man_bus1_range52w(0);
	wire_w_lg_w_man_or2_range84w88w(0) <= wire_w_man_or2_range84w(0) OR wire_w_man_bus2_range86w(0);
	wire_w_lg_w_man_or2_range81w85w(0) <= wire_w_man_or2_range81w(0) OR wire_w_man_bus2_range83w(0);
	wire_w_lg_w_man_or2_range111w115w(0) <= wire_w_man_or2_range111w(0) OR wire_w_man_bus2_range113w(0);
	wire_w_lg_w_man_or2_range108w112w(0) <= wire_w_man_or2_range108w(0) OR wire_w_man_bus2_range110w(0);
	wire_w_lg_w_man_or2_range105w109w(0) <= wire_w_man_or2_range105w(0) OR wire_w_man_bus2_range107w(0);
	wire_w_lg_w_man_or2_range102w106w(0) <= wire_w_man_or2_range102w(0) OR wire_w_man_bus2_range104w(0);
	wire_w_lg_w_man_or2_range99w103w(0) <= wire_w_man_or2_range99w(0) OR wire_w_man_bus2_range101w(0);
	wire_w_lg_w_man_or2_range96w100w(0) <= wire_w_man_or2_range96w(0) OR wire_w_man_bus2_range98w(0);
	wire_w_lg_w_man_or2_range93w97w(0) <= wire_w_man_or2_range93w(0) OR wire_w_man_bus2_range95w(0);
	wire_w_lg_w_man_or2_range90w94w(0) <= wire_w_man_or2_range90w(0) OR wire_w_man_bus2_range92w(0);
	wire_w_lg_w_man_or2_range87w91w(0) <= wire_w_man_or2_range87w(0) OR wire_w_man_bus2_range89w(0);
	wire_w_lg_w_sticky_or_range135w139w(0) <= wire_w_sticky_or_range135w(0) OR wire_w_sticky_bus_range137w(0);
	wire_w_lg_w_sticky_or_range165w169w(0) <= wire_w_sticky_or_range165w(0) OR wire_w_sticky_bus_range167w(0);
	wire_w_lg_w_sticky_or_range168w172w(0) <= wire_w_sticky_or_range168w(0) OR wire_w_sticky_bus_range170w(0);
	wire_w_lg_w_sticky_or_range171w175w(0) <= wire_w_sticky_or_range171w(0) OR wire_w_sticky_bus_range173w(0);
	wire_w_lg_w_sticky_or_range174w178w(0) <= wire_w_sticky_or_range174w(0) OR wire_w_sticky_bus_range176w(0);
	wire_w_lg_w_sticky_or_range177w181w(0) <= wire_w_sticky_or_range177w(0) OR wire_w_sticky_bus_range179w(0);
	wire_w_lg_w_sticky_or_range180w184w(0) <= wire_w_sticky_or_range180w(0) OR wire_w_sticky_bus_range182w(0);
	wire_w_lg_w_sticky_or_range183w187w(0) <= wire_w_sticky_or_range183w(0) OR wire_w_sticky_bus_range185w(0);
	wire_w_lg_w_sticky_or_range186w190w(0) <= wire_w_sticky_or_range186w(0) OR wire_w_sticky_bus_range188w(0);
	wire_w_lg_w_sticky_or_range189w193w(0) <= wire_w_sticky_or_range189w(0) OR wire_w_sticky_bus_range191w(0);
	wire_w_lg_w_sticky_or_range192w196w(0) <= wire_w_sticky_or_range192w(0) OR wire_w_sticky_bus_range194w(0);
	wire_w_lg_w_sticky_or_range138w142w(0) <= wire_w_sticky_or_range138w(0) OR wire_w_sticky_bus_range140w(0);
	wire_w_lg_w_sticky_or_range195w199w(0) <= wire_w_sticky_or_range195w(0) OR wire_w_sticky_bus_range197w(0);
	wire_w_lg_w_sticky_or_range141w145w(0) <= wire_w_sticky_or_range141w(0) OR wire_w_sticky_bus_range143w(0);
	wire_w_lg_w_sticky_or_range144w148w(0) <= wire_w_sticky_or_range144w(0) OR wire_w_sticky_bus_range146w(0);
	wire_w_lg_w_sticky_or_range147w151w(0) <= wire_w_sticky_or_range147w(0) OR wire_w_sticky_bus_range149w(0);
	wire_w_lg_w_sticky_or_range150w154w(0) <= wire_w_sticky_or_range150w(0) OR wire_w_sticky_bus_range152w(0);
	wire_w_lg_w_sticky_or_range153w157w(0) <= wire_w_sticky_or_range153w(0) OR wire_w_sticky_bus_range155w(0);
	wire_w_lg_w_sticky_or_range156w160w(0) <= wire_w_sticky_or_range156w(0) OR wire_w_sticky_bus_range158w(0);
	wire_w_lg_w_sticky_or_range159w163w(0) <= wire_w_sticky_or_range159w(0) OR wire_w_sticky_bus_range161w(0);
	wire_w_lg_w_sticky_or_range162w166w(0) <= wire_w_sticky_or_range162w(0) OR wire_w_sticky_bus_range164w(0);
	aclr <= '0';
	add_1_cout_w <= ((wire_add_sub7_cout AND add_1_w) AND wire_sign_input_reg3_w_lg_q224w(0));
	add_1_w <= (wire_w_lg_w_lg_w_lg_guard_bit_w201w202w203w(0) OR (guard_bit_w AND round_bit_w));
	all_zeroes_w <= ( "0" & "0000000000000000000000000000000");
	barrel_mantissa_input <= ( barrel_zero_padding_w & implied_mantissa_input);
	barrel_zero_padding_w <= (OTHERS => '0');
	below_limit_exceeders <= (((denormal_input_w OR zero_input_w) OR lower_limit_selector) OR nan_input_w);
	below_limit_integer <= (wire_w_lg_w_lg_below_limit_exceeders267w268w OR wire_w_lg_below_limit_exceeders266w);
	below_lower_limit1_w <= wire_cmpr2_aeb;
	below_lower_limit2_w <= wire_cmpr3_alb;
	bias_value_less_1_w <= "01111110";
	bias_value_w <= "01111111";
	clk_en <= '1';
	const_bias_value_add_width_res_w <= "10011110";
	denormal_input_w <= (wire_exp_or_reg4_w_lg_q118w(0) AND man_or_reg4);
	equal_upper_limit_w <= wire_cmpr1_aeb;
	exceed_limit_exceeders <= (wire_w_lg_w_lg_infinity_input_w274w275w(0) AND wire_w_lg_nan_input_w273w(0));
	exceed_limit_integer <= (wire_w_lg_w_lg_exceed_limit_exceeders278w279w OR wire_w_lg_exceed_limit_exceeders277w);
	exceed_upper_limit_w <= wire_cmpr1_agb;
	exp_and <= ( wire_w_lg_w_exp_and_range38w44w & wire_w_lg_w_exp_and_range33w39w & wire_w_lg_w_exp_and_range28w34w & wire_w_lg_w_exp_and_range23w29w & wire_w_lg_w_exp_and_range18w24w & wire_w_lg_w_exp_and_range13w19w & wire_w_lg_w_exp_and_range8w14w & exp_bus(0));
	exp_and_w <= exp_and(7);
	exp_bus <= exponent_input;
	exp_or <= ( wire_w_lg_w_exp_or_range36w42w & wire_w_lg_w_exp_or_range31w37w & wire_w_lg_w_exp_or_range26w32w & wire_w_lg_w_exp_or_range21w27w & wire_w_lg_w_exp_or_range16w22w & wire_w_lg_w_exp_or_range11w17w & wire_w_lg_w_exp_or_range6w12w & exp_bus(0));
	exp_or_w <= exp_or(7);
	exponent_input <= dataa_reg(30 DOWNTO 23);
	guard_bit_w <= wire_altbarrel_shift6_result(23);
	implied_mantissa_input <= ( "1" & mantissa_input_reg);
	infinity_input_w <= (exp_and_reg4 AND wire_man_or_reg4_w_lg_q120w(0));
	infinity_value_w <= (wire_w_lg_w_lg_sign_input_w238w271w OR wire_w_lg_sign_input_w270w);
	int_or1_w <= man_or2(0);
	int_or2_w <= man_or1(0);
	integer_output <= ( sign_input_w & integer_tmp_output);
	integer_post_round <= wire_add_sub7_result;
	integer_pre_round <= lbarrel_shift_w;
	integer_result <= exceed_limit_integer;
	integer_rounded <= (wire_w_lg_w_lg_lowest_integer_selector213w214w OR wire_w_lg_lowest_integer_selector212w);
	integer_rounded_tmp <= (wire_w_lg_w_lg_add_1_w206w207w OR wire_w_lg_add_1_w205w);
	integer_tmp_output <= (wire_w_lg_w_lg_sign_input_w238w239w OR wire_w_lg_sign_input_w237w);
	inv_add_1_adder1_w <= wire_add_sub8_result;
	inv_add_1_adder2_w <= (wire_add_sub8_w_lg_w_lg_cout233w234w OR wire_add_sub8_w_lg_cout232w);
	inv_integer <= (NOT integer_rounded_reg);
	lbarrel_shift_result_w <= wire_altbarrel_shift6_result;
	lbarrel_shift_w <= lbarrel_shift_result_w(53 DOWNTO 23);
	lower_limit_selector <= ((wire_below_lower_limit2_reg4_w_lg_q260w(0) AND wire_w_lg_denormal_input_w258w(0)) AND wire_lowest_int_sel_reg_w_lg_q257w(0));
	lowest_integer_selector <= (below_lower_limit1_reg3 AND man_or_reg3);
	lowest_integer_value <= ( barrel_zero_padding_w & "1");
	man_bus1 <= mantissa_input(10 DOWNTO 0);
	man_bus2 <= mantissa_input(22 DOWNTO 11);
	man_or1 <= ( man_bus1(10) & wire_w_lg_w_man_or1_range47w51w & wire_w_lg_w_man_or1_range50w54w & wire_w_lg_w_man_or1_range53w57w & wire_w_lg_w_man_or1_range56w60w & wire_w_lg_w_man_or1_range59w63w & wire_w_lg_w_man_or1_range62w66w & wire_w_lg_w_man_or1_range65w69w & wire_w_lg_w_man_or1_range68w72w & wire_w_lg_w_man_or1_range71w75w & wire_w_lg_w_man_or1_range74w78w);
	man_or1_w <= man_or1(0);
	man_or2 <= ( man_bus2(11) & wire_w_lg_w_man_or2_range81w85w & wire_w_lg_w_man_or2_range84w88w & wire_w_lg_w_man_or2_range87w91w & wire_w_lg_w_man_or2_range90w94w & wire_w_lg_w_man_or2_range93w97w & wire_w_lg_w_man_or2_range96w100w & wire_w_lg_w_man_or2_range99w103w & wire_w_lg_w_man_or2_range102w106w & wire_w_lg_w_man_or2_range105w109w & wire_w_lg_w_man_or2_range108w112w & wire_w_lg_w_man_or2_range111w115w);
	man_or2_w <= man_or2(0);
	man_or_w <= (man_or1_reg1 OR man_or2_reg1);
	mantissa_input <= dataa_reg(22 DOWNTO 0);
	max_shift_reg_w <= max_shift_reg;
	max_shift_w <= "011110";
	more_than_max_shift_w <= ((max_shift_reg_w AND add_1_cout_w) AND wire_below_lower_limit2_reg3_w_lg_q229w(0));
	nan_input_w <= (exp_and_reg4 AND man_or_reg4);
	neg_infi_w <= ( "1" & "0000000000000000000000000000000");
	padded_exponent_input <= exponent_input;
	pos_infi_w <= ( "0" & "1111111111111111111111111111111");
	power2_value_w <= wire_add_sub4_result(5 DOWNTO 0);
	result <= result_w;
	result_w <= integer_result_reg;
	round_bit_w <= wire_altbarrel_shift6_result(22);
	sign_input <= dataa_reg(31);
	sign_input_w <= sign_input_reg4;
	signed_integer <= ( inv_add_1_adder2_w & inv_add_1_adder1_w);
	sticky_bit_w <= sticky_or(21);
	sticky_bus <= wire_altbarrel_shift6_result(21 DOWNTO 0);
	sticky_or <= ( wire_w_lg_w_sticky_or_range195w199w & wire_w_lg_w_sticky_or_range192w196w & wire_w_lg_w_sticky_or_range189w193w & wire_w_lg_w_sticky_or_range186w190w & wire_w_lg_w_sticky_or_range183w187w & wire_w_lg_w_sticky_or_range180w184w & wire_w_lg_w_sticky_or_range177w181w & wire_w_lg_w_sticky_or_range174w178w & wire_w_lg_w_sticky_or_range171w175w & wire_w_lg_w_sticky_or_range168w172w & wire_w_lg_w_sticky_or_range165w169w & wire_w_lg_w_sticky_or_range162w166w & wire_w_lg_w_sticky_or_range159w163w & wire_w_lg_w_sticky_or_range156w160w & wire_w_lg_w_sticky_or_range153w157w & wire_w_lg_w_sticky_or_range150w154w & wire_w_lg_w_sticky_or_range147w151w & wire_w_lg_w_sticky_or_range144w148w & wire_w_lg_w_sticky_or_range141w145w & wire_w_lg_w_sticky_or_range138w142w & wire_w_lg_w_sticky_or_range135w139w & sticky_bus(0));
	unsigned_integer <= integer_rounded_reg;
	upper_limit_w <= ((wire_sign_input_reg3_w_lg_q224w(0) AND (exceed_upper_limit_reg3 OR equal_upper_limit_reg3)) OR wire_sign_input_reg3_w_lg_q222w(0));
	zero_input_w <= (wire_exp_or_reg4_w_lg_q118w(0) AND wire_man_or_reg4_w_lg_q120w(0));
	wire_w_exp_and_range8w(0) <= exp_and(0);
	wire_w_exp_and_range13w(0) <= exp_and(1);
	wire_w_exp_and_range18w(0) <= exp_and(2);
	wire_w_exp_and_range23w(0) <= exp_and(3);
	wire_w_exp_and_range28w(0) <= exp_and(4);
	wire_w_exp_and_range33w(0) <= exp_and(5);
	wire_w_exp_and_range38w(0) <= exp_and(6);
	wire_w_exp_bus_range10w(0) <= exp_bus(1);
	wire_w_exp_bus_range15w(0) <= exp_bus(2);
	wire_w_exp_bus_range20w(0) <= exp_bus(3);
	wire_w_exp_bus_range25w(0) <= exp_bus(4);
	wire_w_exp_bus_range30w(0) <= exp_bus(5);
	wire_w_exp_bus_range35w(0) <= exp_bus(6);
	wire_w_exp_bus_range40w(0) <= exp_bus(7);
	wire_w_exp_or_range6w(0) <= exp_or(0);
	wire_w_exp_or_range11w(0) <= exp_or(1);
	wire_w_exp_or_range16w(0) <= exp_or(2);
	wire_w_exp_or_range21w(0) <= exp_or(3);
	wire_w_exp_or_range26w(0) <= exp_or(4);
	wire_w_exp_or_range31w(0) <= exp_or(5);
	wire_w_exp_or_range36w(0) <= exp_or(6);
	wire_w_inv_integer_range218w <= inv_integer(30 DOWNTO 15);
	wire_w_man_bus1_range76w(0) <= man_bus1(0);
	wire_w_man_bus1_range73w(0) <= man_bus1(1);
	wire_w_man_bus1_range70w(0) <= man_bus1(2);
	wire_w_man_bus1_range67w(0) <= man_bus1(3);
	wire_w_man_bus1_range64w(0) <= man_bus1(4);
	wire_w_man_bus1_range61w(0) <= man_bus1(5);
	wire_w_man_bus1_range58w(0) <= man_bus1(6);
	wire_w_man_bus1_range55w(0) <= man_bus1(7);
	wire_w_man_bus1_range52w(0) <= man_bus1(8);
	wire_w_man_bus1_range49w(0) <= man_bus1(9);
	wire_w_man_bus2_range113w(0) <= man_bus2(0);
	wire_w_man_bus2_range83w(0) <= man_bus2(10);
	wire_w_man_bus2_range110w(0) <= man_bus2(1);
	wire_w_man_bus2_range107w(0) <= man_bus2(2);
	wire_w_man_bus2_range104w(0) <= man_bus2(3);
	wire_w_man_bus2_range101w(0) <= man_bus2(4);
	wire_w_man_bus2_range98w(0) <= man_bus2(5);
	wire_w_man_bus2_range95w(0) <= man_bus2(6);
	wire_w_man_bus2_range92w(0) <= man_bus2(7);
	wire_w_man_bus2_range89w(0) <= man_bus2(8);
	wire_w_man_bus2_range86w(0) <= man_bus2(9);
	wire_w_man_or1_range47w(0) <= man_or1(10);
	wire_w_man_or1_range74w(0) <= man_or1(1);
	wire_w_man_or1_range71w(0) <= man_or1(2);
	wire_w_man_or1_range68w(0) <= man_or1(3);
	wire_w_man_or1_range65w(0) <= man_or1(4);
	wire_w_man_or1_range62w(0) <= man_or1(5);
	wire_w_man_or1_range59w(0) <= man_or1(6);
	wire_w_man_or1_range56w(0) <= man_or1(7);
	wire_w_man_or1_range53w(0) <= man_or1(8);
	wire_w_man_or1_range50w(0) <= man_or1(9);
	wire_w_man_or2_range84w(0) <= man_or2(10);
	wire_w_man_or2_range81w(0) <= man_or2(11);
	wire_w_man_or2_range111w(0) <= man_or2(1);
	wire_w_man_or2_range108w(0) <= man_or2(2);
	wire_w_man_or2_range105w(0) <= man_or2(3);
	wire_w_man_or2_range102w(0) <= man_or2(4);
	wire_w_man_or2_range99w(0) <= man_or2(5);
	wire_w_man_or2_range96w(0) <= man_or2(6);
	wire_w_man_or2_range93w(0) <= man_or2(7);
	wire_w_man_or2_range90w(0) <= man_or2(8);
	wire_w_man_or2_range87w(0) <= man_or2(9);
	wire_w_sticky_bus_range164w(0) <= sticky_bus(10);
	wire_w_sticky_bus_range167w(0) <= sticky_bus(11);
	wire_w_sticky_bus_range170w(0) <= sticky_bus(12);
	wire_w_sticky_bus_range173w(0) <= sticky_bus(13);
	wire_w_sticky_bus_range176w(0) <= sticky_bus(14);
	wire_w_sticky_bus_range179w(0) <= sticky_bus(15);
	wire_w_sticky_bus_range182w(0) <= sticky_bus(16);
	wire_w_sticky_bus_range185w(0) <= sticky_bus(17);
	wire_w_sticky_bus_range188w(0) <= sticky_bus(18);
	wire_w_sticky_bus_range191w(0) <= sticky_bus(19);
	wire_w_sticky_bus_range137w(0) <= sticky_bus(1);
	wire_w_sticky_bus_range194w(0) <= sticky_bus(20);
	wire_w_sticky_bus_range197w(0) <= sticky_bus(21);
	wire_w_sticky_bus_range140w(0) <= sticky_bus(2);
	wire_w_sticky_bus_range143w(0) <= sticky_bus(3);
	wire_w_sticky_bus_range146w(0) <= sticky_bus(4);
	wire_w_sticky_bus_range149w(0) <= sticky_bus(5);
	wire_w_sticky_bus_range152w(0) <= sticky_bus(6);
	wire_w_sticky_bus_range155w(0) <= sticky_bus(7);
	wire_w_sticky_bus_range158w(0) <= sticky_bus(8);
	wire_w_sticky_bus_range161w(0) <= sticky_bus(9);
	wire_w_sticky_or_range135w(0) <= sticky_or(0);
	wire_w_sticky_or_range165w(0) <= sticky_or(10);
	wire_w_sticky_or_range168w(0) <= sticky_or(11);
	wire_w_sticky_or_range171w(0) <= sticky_or(12);
	wire_w_sticky_or_range174w(0) <= sticky_or(13);
	wire_w_sticky_or_range177w(0) <= sticky_or(14);
	wire_w_sticky_or_range180w(0) <= sticky_or(15);
	wire_w_sticky_or_range183w(0) <= sticky_or(16);
	wire_w_sticky_or_range186w(0) <= sticky_or(17);
	wire_w_sticky_or_range189w(0) <= sticky_or(18);
	wire_w_sticky_or_range192w(0) <= sticky_or(19);
	wire_w_sticky_or_range138w(0) <= sticky_or(1);
	wire_w_sticky_or_range195w(0) <= sticky_or(20);
	wire_w_sticky_or_range141w(0) <= sticky_or(2);
	wire_w_sticky_or_range144w(0) <= sticky_or(3);
	wire_w_sticky_or_range147w(0) <= sticky_or(4);
	wire_w_sticky_or_range150w(0) <= sticky_or(5);
	wire_w_sticky_or_range153w(0) <= sticky_or(6);
	wire_w_sticky_or_range156w(0) <= sticky_or(7);
	wire_w_sticky_or_range159w(0) <= sticky_or(8);
	wire_w_sticky_or_range162w(0) <= sticky_or(9);
	altbarrel_shift6 :  altfp_convert1_altbarrel_shift_grf
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => barrel_mantissa_input,
		distance => power2_value_reg,
		result => wire_altbarrel_shift6_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN added_power2_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN added_power2_reg <= wire_add_sub5_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit1_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit1_reg1 <= below_lower_limit1_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit1_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit1_reg2 <= below_lower_limit1_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit1_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit1_reg3 <= below_lower_limit1_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit2_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit2_reg1 <= below_lower_limit2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit2_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit2_reg2 <= below_lower_limit2_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit2_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit2_reg3 <= below_lower_limit2_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_below_lower_limit2_reg3_w_lg_q229w(0) <= NOT below_lower_limit2_reg3;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit2_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit2_reg4 <= below_lower_limit2_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_below_lower_limit2_reg4_w_lg_q260w(0) <= below_lower_limit2_reg4 AND wire_w_lg_zero_input_w259w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dataa_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dataa_reg <= dataa;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN equal_upper_limit_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN equal_upper_limit_reg1 <= equal_upper_limit_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN equal_upper_limit_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN equal_upper_limit_reg2 <= equal_upper_limit_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN equal_upper_limit_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN equal_upper_limit_reg3 <= equal_upper_limit_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_equal_upper_limit_reg3_w_lg_q220w(0) <= equal_upper_limit_reg3 AND wire_int_or_reg3_w_lg_q219w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg1 <= exceed_upper_limit_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg2 <= exceed_upper_limit_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg3 <= exceed_upper_limit_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_exceed_upper_limit_reg3_w_lg_q221w(0) <= exceed_upper_limit_reg3 OR wire_equal_upper_limit_reg3_w_lg_q220w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg4 <= upper_limit_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg1 <= exp_and_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg2 <= exp_and_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg3 <= exp_and_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg4 <= exp_and_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg1 <= exp_or_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg2 <= exp_or_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg3 <= exp_or_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg4 <= exp_or_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_exp_or_reg4_w_lg_q118w(0) <= NOT exp_or_reg4;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or1_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or1_reg1 <= int_or1_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or2_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or2_reg1 <= int_or2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or_reg2 <= (int_or1_reg1 OR int_or2_reg1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or_reg3 <= int_or_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_int_or_reg3_w_lg_q219w(0) <= int_or_reg3 OR add_1_w;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN integer_result_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN integer_result_reg <= integer_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN integer_rounded_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN integer_rounded_reg <= integer_rounded;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lowest_int_sel_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lowest_int_sel_reg <= lowest_integer_selector;
			END IF;
		END IF;
	END PROCESS;
	wire_lowest_int_sel_reg_w_lg_q257w(0) <= NOT lowest_int_sel_reg;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or1_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or1_reg1 <= man_or1_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or2_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or2_reg1 <= man_or2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or_reg2 <= man_or_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or_reg3 <= man_or_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or_reg4 <= man_or_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_man_or_reg4_w_lg_q120w(0) <= NOT man_or_reg4;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissa_input_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissa_input_reg <= mantissa_input;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN max_shift_exceeder_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN max_shift_exceeder_reg <= more_than_max_shift_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN max_shift_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN max_shift_reg <= wire_max_shift_compare_agb;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN power2_value_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN power2_value_reg <= power2_value_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg1 <= sign_input;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg2 <= sign_input_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg3 <= sign_input_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_sign_input_reg3_w_lg_q222w(0) <= sign_input_reg3 AND wire_exceed_upper_limit_reg3_w_lg_q221w(0);
	wire_sign_input_reg3_w_lg_q224w(0) <= NOT sign_input_reg3;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg4 <= sign_input_reg3;
			END IF;
		END IF;
	END PROCESS;
	add_sub4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_WIDTH => 8,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => exponent_input,
		datab => bias_value_w,
		result => wire_add_sub4_result
	  );
	wire_add_sub5_datab <= "000001";
	add_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 6,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => power2_value_reg,
		datab => wire_add_sub5_datab,
		result => wire_add_sub5_result
	  );
	wire_add_sub7_datab <= "0000000000000000000000000000001";
	add_sub7 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 31,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_sub7_cout,
		dataa => integer_pre_round,
		datab => wire_add_sub7_datab,
		result => wire_add_sub7_result
	  );
	loop42 : FOR i IN 0 TO 15 GENERATE 
		wire_add_sub8_w_lg_w_lg_cout233w234w(i) <= wire_add_sub8_w_lg_cout233w(0) AND wire_w_inv_integer_range218w(i);
	END GENERATE loop42;
	loop43 : FOR i IN 0 TO 15 GENERATE 
		wire_add_sub8_w_lg_cout232w(i) <= wire_add_sub8_cout AND wire_add_sub9_result(i);
	END GENERATE loop43;
	wire_add_sub8_w_lg_cout233w(0) <= NOT wire_add_sub8_cout;
	wire_add_sub8_datab <= "000000000000001";
	add_sub8 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 15,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_sub8_cout,
		dataa => inv_integer(14 DOWNTO 0),
		datab => wire_add_sub8_datab,
		result => wire_add_sub8_result
	  );
	wire_add_sub9_datab <= "0000000000000001";
	add_sub9 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 16,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => inv_integer(30 DOWNTO 15),
		datab => wire_add_sub9_datab,
		result => wire_add_sub9_result
	  );
	cmpr1 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aeb => wire_cmpr1_aeb,
		agb => wire_cmpr1_agb,
		dataa => padded_exponent_input,
		datab => const_bias_value_add_width_res_w
	  );
	cmpr2 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aeb => wire_cmpr2_aeb,
		dataa => exponent_input,
		datab => bias_value_less_1_w
	  );
	cmpr3 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		alb => wire_cmpr3_alb,
		dataa => exponent_input,
		datab => bias_value_w
	  );
	max_shift_compare :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		agb => wire_max_shift_compare_agb,
		dataa => added_power2_reg,
		datab => max_shift_w
	  );

 END RTL; --altfp_convert1_altfp_convert_3tm
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altfp_convert1 IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END altfp_convert1;


ARCHITECTURE RTL OF altfp_convert1 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT altfp_convert1_altfp_convert_3tm
	PORT (
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	altfp_convert1_altfp_convert_3tm_component : altfp_convert1_altfp_convert_3tm
	PORT MAP (
		clock => clock,
		dataa => dataa,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_convert"
-- Retrieval info: CONSTANT: OPERATION STRING "FLOAT2INT"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_DATA NUMERIC "32"
-- Retrieval info: CONSTANT: WIDTH_EXP_INPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_EXP_OUTPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_INT NUMERIC "32"
-- Retrieval info: CONSTANT: WIDTH_MAN_INPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_MAN_OUTPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "32"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: dataa 0 0 32 0 INPUT NODEFVAL "dataa[31..0]"
-- Retrieval info: CONNECT: @dataa 0 0 32 0 dataa 0 0 32 0
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert1.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert1.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert1.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert1_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert1.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert1.cmp TRUE TRUE
-- Retrieval info: LIB_FILE: lpm
