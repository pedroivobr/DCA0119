altfp_convert3_inst : altfp_convert3 PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
