library verilog;
use verilog.vl_types.all;
entity timeSelector_vlg_check_tst is
    port(
        saida           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end timeSelector_vlg_check_tst;
