library verilog;
use verilog.vl_types.all;
entity testes_vlg_vec_tst is
end testes_vlg_vec_tst;
